// audio_system_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module audio_system_tb (
	);

	wire    audio_system_inst_clk_bfm_clk_clk;       // audio_system_inst_clk_bfm:clk -> [audio_system_inst:clk_clk, audio_system_inst_reset_bfm:clk]
	wire    audio_system_inst_reset_bfm_reset_reset; // audio_system_inst_reset_bfm:reset -> audio_system_inst:reset_reset_n

	audio_system audio_system_inst (
		.audio_config_i2c_SDAT   (),                                        // audio_config_i2c.SDAT
		.audio_config_i2c_SCLK   (),                                        //                 .SCLK
		.audio_interface_ADCDAT  (),                                        //  audio_interface.ADCDAT
		.audio_interface_ADCLRCK (),                                        //                 .ADCLRCK
		.audio_interface_BCLK    (),                                        //                 .BCLK
		.audio_interface_DACDAT  (),                                        //                 .DACDAT
		.audio_interface_DACLRCK (),                                        //                 .DACLRCK
		.clk_clk                 (audio_system_inst_clk_bfm_clk_clk),       //              clk.clk
		.key_external_export     (),                                        //     key_external.export
		.led_external_export     (),                                        //     led_external.export
		.reset_reset_n           (audio_system_inst_reset_bfm_reset_reset), //            reset.reset_n
		.switch_external_export  ()                                         //  switch_external.export
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) audio_system_inst_clk_bfm (
		.clk (audio_system_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) audio_system_inst_reset_bfm (
		.reset (audio_system_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (audio_system_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
